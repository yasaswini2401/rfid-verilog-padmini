`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 25.08.2022 10:34:57
// Design Name: 
// Module Name: rx_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// module rx (reset, clk, demodin, bitout, bitclk, rx_overflow_reset, trcal,
//rngbitout);
//////////////////////////////////////////////////////////////////////////////////
module rx_tb();
    reg reset, clk, demodin;
    wire bitout, bitclk, rx_overflow_reset, rngbitout;
    wire [9:0] count;
    wire [9:0] trcal;
    
    reg [1800:0] bitall;
    integer k = 0;
    
    rx r1(.reset(reset),.clk(clk),.demodin(demodin),.bitout(bitout),.bitclk(bitclk),
          .rx_overflow_reset(rx_overflow_reset),.rngbitout(rngbitout),.trcal(trcal), .count(count));
          
    initial begin
        reset = 1;
        clk = 0;
        demodin = 1;
        #0.1
        reset = 0;

        end
    
    always #0.01 clk = ~clk; //2.5MHz clock frequency, bit rate

    initial begin
       bitall = 1801'b1111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111100000000000000000000000011111111111111111111111;
    end


    always@(posedge clk && !reset) begin
    //initial
    
        bitall <= bitall >> 1;
        demodin = bitall;
    end


endmodule